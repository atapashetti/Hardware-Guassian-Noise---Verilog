`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/21/2016 05:11:12 PM
// Design Name: 
// Module Name: cos_sine_TB
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module cos_sine_TB( );

reg clk, rst;
reg [15:0] U1;
wire [15:0] g0, g1;


cos_sine cos_sine1(.clk(clk), 
                   .rst(rst), 
                   .U1(U1), 
                   .g0(g0), 
                   .g1(g1)
                    );
                    
always #10 clk = !clk;

initial begin

	clk = 1'b0;
	rst = 1'b1;

	#30; rst = 1'b0;
	#20; U1 = 16'b0000_0000_0000_0000;
	#20; U1 = 16'b0000_1000_1100_0000;
	#20; U1 = 16'b0011_1111_1111_1110;
	#20; U1 = 16'b0000_0000_0110_1110;

	#20; U1 = 16'b0100_0000_0000_0000;
	#20; U1 = 16'b0100_1000_1100_0000;
	#20; U1 = 16'b0111_1111_1111_1110;
	#20; U1 = 16'b0100_0000_0110_1110;

	#20; U1 = 16'b1000_0000_0000_0000;
	#20; U1 = 16'b1000_1000_1100_0000;
	#20; U1 = 16'b1011_1111_1111_1110;
	#20; U1 = 16'b1000_0000_0110_1110;

	#20; U1 = 16'b1100_0000_0000_0000;
	#20; U1 = 16'b1100_1000_1100_0000;
	#20; U1 = 16'b1111_1111_1111_1110;
	#20; U1 = 16'b1100_0000_0110_1110;

end
endmodule
